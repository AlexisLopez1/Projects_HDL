module mux_nx1(in, select, out);
	parameter SEL = 2;
	parameter DW = 2;
	input data_sel in;
	input logic[SEL-1:0] select;
	output logic[DW-1:0] out;
	
	
	
endmodule 