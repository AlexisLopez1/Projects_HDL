// Copyright (C) 1991-2010 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 10.0 Build 262 08/18/2010 Service Pack 1 SJ Web Edition
// Created on Sat Feb 26 07:12:53 2011

// synthesis message_off 10175

`timescale 1ns/1ns

module FSM_E6 (
    clock,reset,A,B,
    Z);

    input clock;
    input reset;
    input A;
    input B;
    tri0 reset;
    tri0 A;
    tri0 B;
    output Z;
    reg Z;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter S0=0,S1=1,S2=2,S3=3;

    always @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= S0;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or A or B)
    begin
        Z <= 1'b0;
        case (fstate)
            S0: begin
                if ((A == 1'b1))
                    reg_fstate <= S1;
                else if ((A == 1'b0))
                    reg_fstate <= S2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S0;
            end
            S1: begin
                if ((A == 1'b0))
                    reg_fstate <= S0;
                else if ((A == 1'b1))
                    reg_fstate <= S3;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S1;
            end
            S2: begin
                if ((A == 1'b0))
                    reg_fstate <= S2;
                else if ((A == 1'b1))
                    reg_fstate <= S1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S2;

                if ((B == 1'b1))
                    Z <= 1'b1;
                else if ((B == 1'b0))
                    Z <= 1'b0;
                // Inserting 'else' block to prevent latch inference
                else
                    Z <= 1'b0;
            end
            S3: begin
                if ((A == 1'b1))
                    reg_fstate <= S3;
                else if ((A == 1'b0))
                    reg_fstate <= S0;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= S3;

                if ((B == 1'b1))
                    Z <= 1'b1;
                else if ((B == 1'b0))
                    Z <= 1'b0;
                // Inserting 'else' block to prevent latch inference
                else
                    Z <= 1'b0;
            end
            default: begin
                Z <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // Example FSM editor
